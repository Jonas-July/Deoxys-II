package TestIfc;

interface TestIfc;
	method Bool getTestResult();
endinterface

endpackage